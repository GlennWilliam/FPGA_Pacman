module maze (x, y, r, g, b);

	input logic [9:0] x;
	input logic [8:0] y;
	output logic [7:0] r, g, b;
	
	always_comb begin
	
	    // Default color
        r = 0;
        g = 0;
        b = 0;
        
		if(y == 0 || y == 1 || y == 2 || y == 3 || y == 4 || y == 5 ||
		y == 66 || y == 67 || y == 68 || y == 69 || y == 70 || y == 71) begin
		    r <= 0;
		    g <= 0;
		    b <= 255;
		end
		
		else if(x == 0 || x == 1 || x == 2 || x == 3 || x == 4 || x == 5 ||
		x == 90 || x == 91 || x == 92 || x == 93 || x == 94 || x == 95) begin
		    r <= 0;
		    g <= 0;
		    b <= 255;
		end
		
		// 1
		else if (y >= 9 && y <= 11 && x >= 9 && x <= 20 || y >= 9 && y <= 11 && x >= 24 && x <= 71 ||
		y >= 9 && y <= 11 && x >= 75 && x <= 86) begin
		    r <= 0;
		    g <= 0;
		    b <= 255;
		end
		
        else if (y >= 60 && y <= 62 && x >= 9 && x <= 20 || y >= 60 && y <= 62 && x >= 24 && x <= 71 ||
		y >= 60 && y <= 62 && x >= 75 && x <= 86) begin
		    r <= 0;
		    g <= 0;
		    b <= 255;
		end
		
		// 2
		else if (y >= 12 && y <= 14 && x >= 42 && x <= 50) begin
		    r <= 0;
		    g <= 0;
		    b <= 255;
		end
		
		else if (y >= 57 && y <= 59 && x >= 42 && x <= 50) begin
		    r <= 0;
		    g <= 0;
		    b <= 255;
		end
		
		// 3
		else if (y >= 15 && y <= 17 && x >= 9 && x <= 20 || y >= 15 && y <= 17 && x >= 24 && x <= 38 ||
		y >= 15 && y <= 17 && x >= 42 && x <= 50 || y >= 15 && y <= 17 && x >= 54 && x <= 71 ||
		y >= 15 && y <= 17 && x >= 75 && x <= 86) begin
		    r <= 0;
		    g <= 0;
		    b <= 255;
		end
		
		else if (y >= 54 && y <= 56 && x >= 9 && x <= 20 || y >= 54 && y <= 56 && x >= 24 && x <= 38 ||
		y >= 54 && y <= 56 && x >= 42 && x <= 50 || y >= 54 && y <= 56 && x >= 54 && x <= 71 ||
		y >= 54 && y <= 56 && x >= 75 && x <= 86) begin
		    r <= 0;
		    g <= 0;
		    b <= 255;
		end
		
		// 4
		else if (y >= 18 && y <= 20 && x >= 24 && x <= 38 || y >= 18 && y <= 20 && x >= 42 && x <= 50 ||
		y >= 18 && y <= 20 && x >= 54 && x <= 71) begin
		    r <= 0;
		    g <= 0;
		    b <= 255;
		end
		
		else if (y >= 51 && y <= 53 && x >= 24 && x <= 38 || y >= 51 && y <= 53 && x >= 42 && x <= 50 ||
		y >= 51 && y <= 53 && x >= 54 && x <= 71) begin
		    r <= 0;
		    g <= 0;
		    b <= 255;
		end
		
		// 5
		else if (y >= 21 && y <= 26 && x >= 9 && x <= 20 || y >= 21 && y <= 26 && x >= 24 && x <= 38 ||
	    y >= 21 && y <= 26 && x >= 42 && x <= 50 || y >= 21 && y <= 26 && x >= 54 && x <= 71 ||
		y >= 21 && y <= 26 && x >= 75 && x <= 86) begin
		    r <= 0;
		    g <= 0;
		    b <= 255;
		end
		
		else if (y >= 42 && y <= 50 && x >= 9 && x <= 20 || y >= 42 && y <= 50 && x >= 24 && x <= 38 ||
	    y >= 42 && y <= 50 && x >= 42 && x <= 50 || y >= 42 && y <= 50 && x >= 54 && x <= 71 ||
		y >= 42 && y <= 50 && x >= 75 && x <= 86) begin
		    r <= 0;
		    g <= 0;
		    b <= 255;
		end
		
		// 6
		else if (y >= 27 && y <= 29 && x >= 9 && x <= 20 || y >= 27 && y <= 29 && x >= 75 && x <= 86) begin
		    r <= 0;
		    g <= 0;
		    b <= 255;
		end
		
		else if (y >= 39 && y <= 41 && x >= 9 && x <= 20 || y >= 39 && y <= 41 && x >= 75 && x <= 86) begin
		    r <= 0;
		    g <= 0;
		    b <= 255;
		end
		
		else if (y >= 30 && y <= 38 && x >= 9 && x <= 20 || y >= 30 && y <= 38 && x >= 24 && x <= 71 ||
		y >= 30 && y <= 38 && x >= 75 && x <= 86) begin
		    r <= 0;
		    g <= 0;
		    b <= 255;
		end
	
	end
	
endmodule